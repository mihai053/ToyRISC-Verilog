module programmemory(
	input [15:0] instrAddr,
	output reg [31:0] instruction,
	input clock,
	input reset
    );
	 reg [31:0] mem [0:65535];
	 
	 always @(posedge clock)
	 if(reset)
		begin
			instruction<=0;
			//////////////////////////////////////////////////
			///////////////codul lui Claudiu//////////////////
			/*mem[0] =32'b010111_00000_00000_00000_00000000010;
			mem[1] =32'b010111_00001_00000_00000_00000000001;
			mem[2] =32'b010111_00010_00000_00000_00000000100;
			mem[3] =32'b111110_00000_00001_00010_00000000000;
			mem[4] =32'b000111_00011_00000_00000_00000011111;
			mem[31] =32'b000000_00000_00000_00000_00000000000;
			mem[32] =32'b110010_00100_00001_00010_00000000000;
			mem[33] =32'b101000_00000_00000_00010_00000000000;
			mem[34] =32'b000101_00000_00011_00000_00000000000;*/
			//////////////////////////////////////////////////
			////////////////codul lui Tache///////////////////
			mem[0] =32'b010111_00000_00000_00000_00000000101;
			mem[1] =32'b000011_00000_00001_00000_00000011111;
			mem[2] =32'b000111_00101_00000_00000_00000011111;
			mem[3] =32'b000010_00000_00001_00010_00000000101;
			mem[4] =32'b000110_00000_00000_00000_00000000010;
			mem[5] =32'b110010_00001_00001_00000_00000000000;
			mem[6] =32'b110001_00000_00000_00010_00000000000;
			mem[7] =32'b000101_00000_11111_00000_00000000000;
			mem[8] =32'b010111_00000_00011_00000_00000000000;
			//////////////////////////////////////////////////
		end 
	else
		instruction <= mem[instrAddr];   
endmodule
   




